* Only a small resistor 
rm b c 3.16G
vm c 0 dc 0.060
cm b 0 3.1416p
i1 b 0 pulse(0p 10p 0 0.1m 0.1m 0.05 0.1) 

.CONTROL
tran 10m 100ms
plot v(b)
.ENDC

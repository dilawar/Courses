* With 1000 Hz pulse
rm b c 3.16G
vm c 0 dc 0.060
cm b 0 3.1416p
i1 b 0 pulse(0p 10p 0 0.1n 0.1n 0.0005 0.001) 

.CONTROL
set hcopypscolor=1
tran 0.1m 0.1
plot v(b)
hardcopy plot_1000hz.ps v(b)
.ENDC
